*case_2.sp comment
R1 1 2 100
C1 2 0 1p
R2 2 0 100
V1 1 0 DC 1
.DC V1 0 10 1
.PRINT DC V(2)
.PLOT DC V(2)
.END
